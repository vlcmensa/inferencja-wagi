/*
================================================================================
Isolated Testbench for Inference Module
================================================================================

Purpose: Test inference.v in isolation using exact same data preparation as
         Python simulation to eliminate all other error sources.

Strategy:
  1. Load actual weights and biases from .mem files
  2. Load preprocessed test vectors generated by Python
  3. Run inference on each test case
  4. Compare results with expected scores from Python simulation
  5. Report any mismatches

================================================================================
*/

`timescale 1ns / 1ps

module tb_inference_isolated();

    // Parameters
    parameter NUM_PIXELS = 784;
    parameter NUM_CLASSES = 10;
    parameter NUM_TEST_CASES = 100;
    
    // Clock and Reset
    reg clk;
    reg rst;
    
    // Memory Interfaces
    wire [12:0] weight_addr;
    reg  [7:0]  weight_data;
    wire [3:0]  bias_addr;
    reg  [31:0] bias_data;
    wire [9:0]  input_addr;
    reg  [7:0]  input_pixel;
    
    // Control
    reg weights_ready;
    reg start_inference;
    
    // Outputs
    wire [3:0] predicted_digit;
    wire inference_done;
    wire busy;
    
    // Class scores
    wire signed [31:0] class_score_0;
    wire signed [31:0] class_score_1;
    wire signed [31:0] class_score_2;
    wire signed [31:0] class_score_3;
    wire signed [31:0] class_score_4;
    wire signed [31:0] class_score_5;
    wire signed [31:0] class_score_6;
    wire signed [31:0] class_score_7;
    wire signed [31:0] class_score_8;
    wire signed [31:0] class_score_9;
    
    // Test data storage - FLATTENED arrays for proper $readmemh loading
    reg [7:0] weights_mem [0:7839];
    reg [31:0] biases_mem [0:9];
    reg [7:0] test_pixels_flat [0:78399];      // 100 tests * 784 pixels = 78400
    reg signed [31:0] expected_scores_flat [0:999];  // 100 tests * 10 scores = 1000
    reg [3:0] expected_predictions [0:99];
    reg [3:0] true_labels [0:99];
    
    // Test control
    integer test_idx;
    integer pass_count;
    integer fail_count;
    integer j;
    integer file_check;  // For file loading error checking
    reg signed [31:0] max_error;
    reg scores_match;
    reg signed [31:0] fpga_scores [0:9];
    reg signed [31:0] diff;
    
    // Instantiate the Unit Under Test (UUT)
    inference uut (
        .clk(clk),
        .rst(rst),
        .weight_addr(weight_addr),
        .weight_data(weight_data),
        .bias_addr(bias_addr),
        .bias_data(bias_data),
        .weights_ready(weights_ready),
        .start_inference(start_inference),
        .input_pixel(input_pixel),
        .input_addr(input_addr),
        .predicted_digit(predicted_digit),
        .inference_done(inference_done),
        .busy(busy),
        .class_score_0(class_score_0),
        .class_score_1(class_score_1),
        .class_score_2(class_score_2),
        .class_score_3(class_score_3),
        .class_score_4(class_score_4),
        .class_score_5(class_score_5),
        .class_score_6(class_score_6),
        .class_score_7(class_score_7),
        .class_score_8(class_score_8),
        .class_score_9(class_score_9)
    );
    
    // Clock Generation: 100MHz
    always #5 clk = ~clk;
    
    // ========================================================================
    // Memory Interface Logic
    // ========================================================================
    
    // Weight Memory
    always @(posedge clk) begin
        if (weight_addr < 7840)
            weight_data <= weights_mem[weight_addr];
        else
            weight_data <= 8'd0;
    end
    
    // Bias Memory
    always @(posedge clk) begin
        if (bias_addr < 10)
            bias_data <= biases_mem[bias_addr];
        else
            bias_data <= 32'd0;
    end
    
    // Input Pixel Memory (access flattened array)
    always @(posedge clk) begin
        if (input_addr < 784)
            input_pixel <= test_pixels_flat[test_idx * 784 + input_addr];
        else
            input_pixel <= 8'd0;
    end
    
    // ========================================================================
    // Load Memory Files
    // ========================================================================
    initial begin
        $display("================================================================================");
        $display("Loading Memory Files...");
        $display("================================================================================");
        $display("Current working directory for file loading:");
        $display("  (Vivado runs from simulation directory)");
        $display("");
        
        // Load weights with error checking
        file_check = $fopen("../../outputs/mem/W.mem", "r");
        if (file_check == 0) begin
            $display("ERROR: Cannot open ../../outputs/mem/W.mem");
            $display("  Make sure you run from regresja/inference/tb/ directory");
            $finish;
        end
        $fclose(file_check);
        $readmemh("../../outputs/mem/W.mem", weights_mem);
        $display("  [OK] Loaded weights: 7840 entries");
        
        // Load biases with error checking
        file_check = $fopen("../../outputs/mem/B.mem", "r");
        if (file_check == 0) begin
            $display("ERROR: Cannot open ../../outputs/mem/B.mem");
            $finish;
        end
        $fclose(file_check);
        $readmemh("../../outputs/mem/B.mem", biases_mem);
        $display("  [OK] Loaded biases: 10 entries");
        
        // Load test vectors (flattened format) with error checking
        file_check = $fopen("test_vectors_pixels.mem", "r");
        if (file_check == 0) begin
            $display("ERROR: Cannot open test_vectors_pixels.mem");
            $display("  Run generate_test_vectors.py first!");
            $display("  Files must be in same directory as testbench");
            $finish;
        end
        $fclose(file_check);
        $readmemh("test_vectors_pixels.mem", test_pixels_flat);
        $display("  [OK] Loaded pixel vectors: 78400 values");
        
        file_check = $fopen("test_vectors_scores.mem", "r");
        if (file_check == 0) begin
            $display("ERROR: Cannot open test_vectors_scores.mem");
            $finish;
        end
        $fclose(file_check);
        $readmemh("test_vectors_scores.mem", expected_scores_flat);
        $display("  [OK] Loaded score vectors: 1000 values");
        
        file_check = $fopen("test_vectors_meta.mem", "r");
        if (file_check == 0) begin
            $display("ERROR: Cannot open test_vectors_meta.mem");
            $finish;
        end
        $fclose(file_check);
        $readmemh("test_vectors_meta.mem", expected_predictions);
        $display("  [OK] Loaded predictions: 100 values");
        
        file_check = $fopen("test_vectors_labels.mem", "r");
        if (file_check == 0) begin
            $display("ERROR: Cannot open test_vectors_labels.mem");
            $finish;
        end
        $fclose(file_check);
        $readmemh("test_vectors_labels.mem", true_labels);
        $display("  [OK] Loaded labels: 100 values");
        
        $display("  [OK] Loaded test vectors: %0d test cases", NUM_TEST_CASES);
        $display("================================================================================\n");
    end
    
    // ========================================================================
    // Test Sequence
    // ========================================================================
    initial begin
        $display("================================================================================");
        $display("Isolated Testbench for inference.v");
        $display("================================================================================");
        $display("Testing inference.v in complete isolation using:");
        $display("  - Real weight and bias files from training");
        $display("  - Preprocessed test vectors from Python (same as UART sends)");
        $display("  - Expected scores from Python simulation (with overflow)");
        $display("================================================================================\n");
        
        // Initialize
        clk = 0;
        rst = 1;
        weights_ready = 0;
        start_inference = 0;
        test_idx = 0;
        pass_count = 0;
        fail_count = 0;
        
        // Reset
        #100;
        rst = 0;
        #20;
        
        $display("[%0t] Starting Isolated Inference Tests\n", $time);
        weights_ready = 1;
        
        // Run tests on all test cases
        for (test_idx = 0; test_idx < NUM_TEST_CASES; test_idx = test_idx + 1) begin
            $display("================================================================================");
            $display("Test Case %0d / %0d", test_idx + 1, NUM_TEST_CASES);
            $display("================================================================================");
            $display("  True Label:         %0d", true_labels[test_idx]);
            $display("  Expected Pred:      %0d (from Python sim)", expected_predictions[test_idx]);
            
            // Start inference
            #10 start_inference = 1;
            #10 start_inference = 0;
            
            // Wait for completion
            wait(inference_done);
            #20;
            
            // Collect FPGA scores
            fpga_scores[0] = class_score_0;
            fpga_scores[1] = class_score_1;
            fpga_scores[2] = class_score_2;
            fpga_scores[3] = class_score_3;
            fpga_scores[4] = class_score_4;
            fpga_scores[5] = class_score_5;
            fpga_scores[6] = class_score_6;
            fpga_scores[7] = class_score_7;
            fpga_scores[8] = class_score_8;
            fpga_scores[9] = class_score_9;
            
            // Verify results
            $display("  FPGA Pred:          %0d", predicted_digit);
            $display("\n  Score Comparison:");
            $display("  Class | Expected      | FPGA          | Difference");
            $display("  ------|---------------|---------------|---------------");
            
            scores_match = 1;
            max_error = 0;
            
            // Compare all class scores (access flattened array)
            for (j = 0; j < 10; j = j + 1) begin
                diff = fpga_scores[j] - expected_scores_flat[test_idx * 10 + j];
                
                if (fpga_scores[j] !== expected_scores_flat[test_idx * 10 + j]) begin
                    scores_match = 0;
                    if ($signed(diff) < 0) begin
                        if (-diff > max_error) max_error = -diff;
                    end else begin
                        if (diff > max_error) max_error = diff;
                    end
                end
                
                $display("    %0d   | %13d | %13d | %13d %s",
                        j, expected_scores_flat[test_idx * 10 + j], fpga_scores[j], diff,
                        (fpga_scores[j] !== expected_scores_flat[test_idx * 10 + j]) ? "<-- MISMATCH" : "");
            end
            
            // Check overall result
            $display("\n  Max Score Error:    %0d", max_error);
            $display("  Scores Match:       %s", scores_match ? "YES" : "NO");
            $display("  Pred Match:         %s", (predicted_digit == expected_predictions[test_idx]) ? "YES" : "NO");
            
            if (scores_match && (predicted_digit == expected_predictions[test_idx])) begin
                $display("  Result:             PASS");
                pass_count = pass_count + 1;
            end else begin
                $display("  Result:             FAIL");
                fail_count = fail_count + 1;
            end
            
            $display("");
            
            // Small delay between tests
            #50;
        end
        
        // Final Summary
        $display("\n================================================================================");
        $display("FINAL RESULTS");
        $display("================================================================================");
        $display("Total Tests:        %0d", NUM_TEST_CASES);
        $display("Passed:             %0d", pass_count);
        $display("Failed:             %0d", fail_count);
        $display("Pass Rate:          %.1f%%", (pass_count * 100.0) / NUM_TEST_CASES);
        $display("================================================================================");
        
        if (fail_count == 0) begin
            $display("\nALL TESTS PASSED");
            $display("inference.v is computing correctly!");
            $display("The mismatch problem is NOT in inference.v");
            $display("Check other modules: UART, image_loader, weight_loader, etc.");
        end else begin
            $display("\nTESTS FAILED");
            $display("inference.v has computation errors!");
            $display("Review the detailed comparisons above.");
            $display("Possible issues:");
            $display("  - Pipeline timing bug");
            $display("  - Sign extension error");
            $display("  - Accumulator overflow handling");
            $display("  - Weight/bias memory addressing");
        end
        $display("================================================================================\n");
        
        #100;
        $finish;
    end
    
    // Timeout watchdog
    initial begin
        #100000000;  // 100ms timeout
        $display("\nERROR: Simulation timeout!");
        $finish;
    end

endmodule